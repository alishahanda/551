module PID #(parameter fast_sim = 1) (clk, rst_n, vld, rider_off, ptch, ptch_rt, pwr_up, PID_cntrl, ss_tmr);

input clk, rst_n, vld, rider_off, pwr_up;
input [15:0] ptch;
input [15:0] ptch_rt;
output [11:0] PID_cntrl;
output [7:0] ss_tmr;

logic signed [9:0] ptch_err_sat;
logic signed [17:0] ptch_err_sat_sign_ext;
logic signed [17:0] integrator;
logic signed [14:0] P_term;
logic signed [14:0] I_term;
logic signed [12:0] D_term;
logic signed [15:0] PID_cntrl_pre_sat;
logic signed [17:0] accumulator;
logic signed valid, ov;
logic signed [26:0] soft_start_ff;
logic signed [26:0] ss_tmr_incr;
logic signed [14:0] integrator_val_for_I_term;

localparam P_COEFF = 5'h0C;

//generate conditional
generate if (fast_sim) begin
		assign ss_tmr_incr = 27'd256; //If fast_sim, we increment ss_tmr by 256 every clock (instead of by 1 every clk)
		assign integrator_val_for_I_term = (!integrator[17] && |integrator[17:15]) ? 15'h3FFF : 
						((integrator[17] && !(&integrator[17:15])) ? 15'h4000 : 
						integrator[15:1]); //saturation logic
	end else begin
		assign ss_tmr_incr = 27'd1;
		assign integrator_val_for_I_term = {{3{integrator[17]}}, integrator[17:6]};
	end
endgenerate

//forming saturated 10-bit error term
assign ptch_err_sat = (~ptch[15] && |ptch[14:9]) ? 10'h1FF : 
					  ((ptch[15] && ~(&ptch[14:9])) ? 10'h200 : 
					  ptch[9:0]) ; //saturate ptch to 10 bit value
					  
//sign extend ptch_err_sat to 18 bits					  
assign ptch_err_sat_sign_ext = {{8{ptch_err_sat[9]}}, ptch_err_sat};

assign accumulator = ptch_err_sat_sign_ext + integrator;

//check for overflow
//overflow occurs if both inputs are positive and output is negative or vice-versa
assign ov = ((ptch_err_sat_sign_ext[17] && integrator[17] && ~accumulator[17]) || 
			(~ptch_err_sat_sign_ext[17] && ~integrator[17] && accumulator[17]));
assign valid = vld & ~ov;

always_ff@(posedge clk, negedge rst_n) begin
	if (!rst_n) 
		integrator <= 'b0;
	else if (rider_off)
		integrator <= 18'b0;
	else if (valid)
		integrator <= accumulator;
end 

assign P_term = ptch_err_sat * $signed(P_COEFF); //signed multiplication

assign I_term = integrator_val_for_I_term; //I_term generated by generate if block depending on value of fast_sim

//D_term = one's comp of (ptch_rt / 64)
assign D_term = ~({{3{ptch_rt[15]}}, ptch_rt[15:6]}); //divide by 64 is same as ARS by 6

//summing up sign extended P_term, D_term and I_term
assign PID_cntrl_pre_sat = {P_term[14], P_term[14:0]} + {I_term[14], I_term[14:0]} + {{3{D_term[12]}}, D_term[12:0]};

assign PID_cntrl = (~PID_cntrl_pre_sat[15] && |PID_cntrl_pre_sat[14:11]) ? 12'h7FF: 
					  ((PID_cntrl_pre_sat[15] && ~(&PID_cntrl_pre_sat[14:11])) ? 12'h800 : 
					  PID_cntrl_pre_sat[11:0]); //saturate to 13 bit value

//Soft start timer
always_ff@(posedge clk, negedge rst_n) begin
	if(!rst_n) 
		soft_start_ff <= 'b0;
	else if (!pwr_up)
		soft_start_ff <= 'h0;
	else if (!(&soft_start_ff[26:8]))
		soft_start_ff <= soft_start_ff + ss_tmr_incr; //incr value determined by generate if block based on value of fast_sim		
end 

assign ss_tmr = soft_start_ff[26:19];

endmodule
